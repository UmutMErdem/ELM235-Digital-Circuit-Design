`timescale 1ns/1ps
module tb_lab3_g7_p5();
logic [3:0] I;
logic [15:0] Q1, Q2;
logic F1, F2;

lab3_g7_p5 dut0(I,Q1,Q2,F1,F2);
initial begin
	I[3]=0; I[2]=0; I[1]=0; I[0]=0; #10
	I[3]=0; I[2]=0; I[1]=0; I[0]=1; #10
	I[3]=0; I[2]=0; I[1]=1; I[0]=0; #10
	I[3]=0; I[2]=0; I[1]=1; I[0]=1; #10
	I[3]=0; I[2]=1; I[1]=0; I[0]=0; #10
	I[3]=0; I[2]=1; I[1]=0; I[0]=1; #10
	I[3]=0; I[2]=1; I[1]=1; I[0]=0; #10
	I[3]=0; I[2]=1; I[1]=1; I[0]=1; #10
	I[3]=1; I[2]=0; I[1]=0; I[0]=0; #10
	I[3]=1; I[2]=0; I[1]=0; I[0]=1; #10
	I[3]=1; I[2]=0; I[1]=1; I[0]=0; #10
	I[3]=1; I[2]=0; I[1]=1; I[0]=1; #10
	I[3]=1; I[2]=1; I[1]=0; I[0]=0; #10
	I[3]=1; I[2]=1; I[1]=0; I[0]=1; #10
	I[3]=1; I[2]=1; I[1]=1; I[0]=0; #10
	I[3]=1; I[2]=1; I[1]=1; I[0]=1; #10
$stop;
end
endmodule
