`timescale 1ns/1ps
module tb_lab3_g7_p4();
logic S;
logic [2:0] I_3;
logic [3:0] I_4;
logic [7:0] Q_8;
logic [15:0] Q_16;

lab3_g7_p4 dut0(S, I_4, Q_16);
decoder4x16 decoder4x16(I_4[3:0], Q_16[15:0]);

initial begin
	I_4[3]=0; I_4[2]=0; I_4[1]=0; I_4[0]=0; #10
	I_4[3]=0; I_4[2]=0; I_4[1]=0; I_4[0]=1; #10
	I_4[3]=0; I_4[2]=0; I_4[1]=1; I_4[0]=0; #10
	I_4[3]=0; I_4[2]=0; I_4[1]=1; I_4[0]=1; #10
	I_4[3]=0; I_4[2]=1; I_4[1]=0; I_4[0]=0; #10
	I_4[3]=0; I_4[2]=1; I_4[1]=0; I_4[0]=1; #10
	I_4[3]=0; I_4[2]=1; I_4[1]=1; I_4[0]=0; #10
	I_4[3]=0; I_4[2]=1; I_4[1]=1; I_4[0]=1; #10
	I_4[3]=1; I_4[2]=0; I_4[1]=0; I_4[0]=0; #10
	I_4[3]=1; I_4[2]=0; I_4[1]=0; I_4[0]=1; #10
	I_4[3]=1; I_4[2]=0; I_4[1]=1; I_4[0]=0; #10
	I_4[3]=1; I_4[2]=0; I_4[1]=1; I_4[0]=1; #10
	I_4[3]=1; I_4[2]=1; I_4[1]=0; I_4[0]=0; #10
	I_4[3]=1; I_4[2]=1; I_4[1]=0; I_4[0]=1; #10
	I_4[3]=1; I_4[2]=1; I_4[1]=1; I_4[0]=0; #10
	I_4[3]=1; I_4[2]=1; I_4[1]=1; I_4[0]=1; #10
	$stop;
end
endmodule
/*
lab3_g7_p4 dut0(S, I_3, Q_8);

decoder3x8 decoder3x8(S, I_3[2:0], Q_8[7:0]);
initial begin
	S=1; I_3[2]=0; I_3[1]=0; I_3[0]=0; #10
	I_3[2]=0; I_3[1]=0; I_3[0]=1; #10
	I_3[2]=0; I_3[1]=1; I_3[0]=0; #10
	I_3[2]=0; I_3[1]=1; I_3[0]=1; #10
	I_3[2]=1; I_3[1]=0; I_3[0]=0; #10
	I_3[2]=1; I_3[1]=0; I_3[0]=1; #10
	I_3[2]=1; I_3[1]=1; I_3[0]=0; #10
	I_3[2]=1; I_3[1]=1; I_3[0]=1; #10
	$stop;
end
endmodule
*/
