`timescale 1ns/1ps
module tb_lab2_g7_p2();
  logic [3:0] x;
  logic [6:0] sev_segments;
  
  lab2_g7_p2 dut0(x, sev_segments);
  
initial begin
 	x[3] = 0; x[2] = 0; x[1] = 0; x[0]=0; 	#10 // 0000
	x[0] = 1;		     	  	#10 // 0001
	x[1] = 1; x[0] = 0;	     	  	#10 // 0010
	x[0] = 1;		     	  	#10 // 0011
	x[2] = 1; x[1] = 0; x[0] = 0; 	  	#10 // 0100
	x[0] = 1;		     	  	#10 // 0101
	x[1] = 1; x[0] = 0;	     	  	#10 // 0110
	x[0] = 1;		     	  	#10 // 0111
	x[3] = 1; x[2] = 0; x[1] = 0; x[0]=0; 	#10 // 1000
	x[0] = 1;		     	  	#10 // 1001
	x[1] = 1; x[0] = 0;	     	  	#10 // 1010
	x[0] = 1;		     	  	#10 // 1011
	x[2] = 1; x[1] = 0; x[0] = 0; 	  	#10 // 1100
	x[0] = 1;		     	  	#10 // 1101
	x[1] = 1; x[0] = 0;	     	  	#10 // 1110
	x[0] = 1;		     	  	#10 // 1111
	$stop;
end
endmodule