`timescale 1ns/1ps
module tb_lab4_g7_p2();
logic [4:0] A, B;
logic Cin;
logic [4:0] S;
logic Cout;

lab4_g7_p2 dut0(A, B, Cin, S, Cout);

initial begin
	A=5'b10001; B=5'b10101; Cin=0; 	#10
	A=5'b10110; B=5'b10000;		#10
	A=5'b10110; B=5'b10111;		#10
	A=5'b01001; B=5'b01011;		#10
	A=5'b01010; B=5'b00110;		#10
	A=5'b01010; B=5'b11111;		#10
	A=5'b01110; B=5'b00110;		#10
	A=5'b10111; B=5'b10110;		#10
	A=5'b01011; B=5'b00001;		#10
	A=5'b01111; B=5'b11110;		#10
	A=5'b11011; B=5'b00111;		#10
	A=5'b10101; B=5'b10111;		#10
	A=5'b10011; B=5'b01100;		#10
	A=5'b11011; B=5'b10110;		#10
	A=5'b01010; B=5'b10111;		#10
	A=5'b00001; B=5'b01000;		#10
	$stop;
end
endmodule
