`timescale 1ns/1ps
module tb_lab2_g7_p1();
  logic A, B, C, D;
  logic X, Y;
  
  lab2_g7_p1 dut0(A, B, C, D, X, Y);
  
initial begin
  	A = 0; B = 0; C = 0; D=0; #10 // 0000
	D = 1;		     	  #10 // 0001
	C = 1; D = 0;	     	  #10 // 0010
	D = 1;		     	  #10 // 0011
	B = 1; C = 0; D = 0; 	  #10 // 0100
	D = 1;		     	  #10 // 0101
	C = 1; D = 0;	     	  #10 // 0110
	D = 1;		     	  #10 // 0111
	A = 1; B = 0; C = 0; D=0; #10 // 1000
	D = 1;		     	  #10 // 1001
	C = 1; D = 0;	     	  #10 // 1010
	D = 1;		     	  #4  // 1011
	C=0;			  #2  // 1011
	C=1;			  #4  // 1011
	B = 1; C = 0; D = 0; 	  #10 // 1100
	D = 1;		     	  #10 // 1101
	C = 1; D = 0;	     	  #10 // 1110
	D = 1;		     	  #10 // 1111
	$stop;
end
endmodule