`timescale 1ns/1ps
module tb_lab4_g7_p3();
logic [31:0] a, b;
logic [3:0] op;
logic [31:0] s;
logic n, z, v, c, hata;

lab4_g7_p3 dut0(a, b, op, s, n, z, v, c, hata);

initial begin
	a=32'h81000003; b=32'h80000007; op=4'b0000; #10
	a=32'h81000003; b=32'h80000007; op=4'b1000; #10
	a=32'h81000003; b=32'h80000007; op=4'b0001; #10
	a=32'h81000003; b=32'h80000007; op=4'b0010; #10
	a=32'h81000003; b=32'h80000007; op=4'b0011; #10
	a=32'h81000003; b=32'h80000007; op=4'b0100; #10
	a=32'h81000003; b=32'h80000007; op=4'b0101; #10
	a=32'h81000003; b=32'h80000007; op=4'b1101; #10
	a=32'h81000003; b=32'h80000007; op=4'b0110; #10
	a=32'h81000003; b=32'h80000007; op=4'b0111; #10
	a=32'h81000003; b=32'h80000007; op=4'b1111; #10
	a=32'h81000003; b=32'h80000007; op=4'b1011; #10
	$stop;
end
endmodule